
module Hamming_Encoder(
    output [7:0] data_out,
    input [3:0] data_in,
    input clk, rstn
    );

// **** TODO **** //



// ************** //

endmodule