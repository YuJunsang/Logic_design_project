
module Hamming_Decoder(
    output [3:0] data_out,
    output err_uncorrectable, err_correctable,
    input [7:0] data_in,
    input clk, rstn
    );

// **** TODO **** //



// ************** //

endmodule
