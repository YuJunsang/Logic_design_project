
module Error_Injection(
        output [7:0] data_out,
        input [7:0] data_in,
        input btn1, btn2,
        input clk, rstn
    );

// **** TODO **** //



// ************** // 

endmodule